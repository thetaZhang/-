module FrequencyMeter (
    input Fxin,
    inout Clk,
    output Frequency
);
    reg[]
endmodule